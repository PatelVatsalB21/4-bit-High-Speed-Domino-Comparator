VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cmp
  CLASS BLOCK ;
  FOREIGN cmp ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.670 BY 34.390 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 35.620 28.890 39.620 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 35.620 17.850 39.620 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END A[3]
  PIN B[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END B[0]
  PIN B[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 24.900 21.800 28.900 22.400 ;
    END
  END B[1]
  PIN B[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END B[2]
  PIN B[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END B[3]
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 15.280 23.000 16.880 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 12.560 23.000 14.160 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 35.620 6.810 39.620 ;
    END
  END clk
  PIN out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 24.900 5.480 28.900 6.080 ;
    END
  END out
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 23.000 27.285 ;
      LAYER met1 ;
        RECT 0.070 26.080 23.670 27.440 ;
        RECT 28.130 26.080 28.450 26.140 ;
        RECT 0.070 25.940 28.450 26.080 ;
        RECT 0.070 10.640 23.670 25.940 ;
        RECT 28.130 25.880 28.450 25.940 ;
      LAYER met2 ;
        RECT 6.600 34.390 6.740 35.620 ;
        RECT 17.640 34.390 17.780 35.620 ;
        RECT 0.100 4.280 23.670 34.390 ;
        RECT 28.680 26.250 28.820 35.620 ;
        RECT 28.220 26.170 28.820 26.250 ;
        RECT 28.160 26.110 28.820 26.170 ;
        RECT 28.160 25.850 28.420 26.110 ;
        RECT 0.650 3.670 10.850 4.280 ;
        RECT 11.690 3.670 21.890 4.280 ;
        RECT 22.730 3.670 23.670 4.280 ;
      LAYER met3 ;
        RECT 4.400 32.280 23.670 33.145 ;
        RECT 4.000 22.250 23.670 32.280 ;
        RECT 4.000 21.950 24.900 22.250 ;
        RECT 4.000 17.360 23.670 21.950 ;
        RECT 4.400 15.960 23.670 17.360 ;
        RECT 4.000 5.930 23.670 15.960 ;
        RECT 4.000 5.630 24.900 5.930 ;
        RECT 4.000 5.615 23.670 5.630 ;
      LAYER met4 ;
        RECT 7.630 10.640 20.885 27.440 ;
      LAYER met5 ;
        RECT 5.520 18.480 23.000 25.040 ;
  END
END cmp
END LIBRARY

